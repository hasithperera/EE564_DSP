----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:48:03 01/07/2016 
-- Design Name: 
-- Module Name:    top - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity top is
    Port ( -- KC705 200 MHz system clock
           SYSCLK_P : in STD_LOGIC; --! KC705 on-board 200 MHz clock generated by a crystal oscillator 
           SYSCLK_N : in STD_LOGIC;

           -- KC705 row of LEDs
		   GPIO_LED: out  STD_LOGIC_VECTOR(7 downto 0); --! Row of 8 leds on the KC705

                    ------------------------------------
            -- KC705 GMII PHY Gigabit Ethernet Interface (Marvell Alaska 10-100-1000BASE-T PHY)
            ------------------------------------
            PHY_RXCLK : in  STD_LOGIC; --! Receive byte clock recovered  by the PHY chip
            PHY_TXER: out STD_LOGIC; --! Enabled to transmit an error condition to the PHY
            PHY_RESET_L: out STD_LOGIC; --! Active LOW PHY reset
            PHY_RXCTRL_RXDV: in  STD_LOGIC; --! RX Data Valid flag from the PHY
            PHY_RXD: in  STD_LOGIC_VECTOR(7 downto 0); -- RX Data from the PHY

            PHY_TXC_GTXCLK: out STD_LOGIC; --! 125 MHz clock provided to the PHY to clock the Tx bus 
            PHY_TXCTL_TXEN: out STD_LOGIC; --! Indicates that valid data is presented on the PHY TX bus.
            PHY_TXD: out  STD_LOGIC_VECTOR(7 downto 0); --! Tx Data bus to the PHY
            PHY_TXCLK: in STD_LOGIC --! 125 MHz TX clock supplied *by* the PHY. This is not used as we generate our own clock internally.
         );



end top;

architecture Behavioral of top is

-- Clocks & global reset
signal CLK125: std_logic; --! 125 MHz clock for the command interface and the Ethernet communications  
signal CLK200: std_logic; --! 200 MHz system clock from the carrier board  
signal CLK200_MMCM_NOBUF : std_logic; --! 200 MHz clock generated by a MMCM, *without* a BUFG. Is meant to be connected to the BUFGMUX that select the antenna processing clock. Cannot clock logic.
signal CLK25: std_logic; -- 25 MHz clock  
signal CORR_CLK: std_logic; --! Correlator clock, derived from the carrier board. 
signal CORR_CLK_MMCM: std_logic; --! Correlator clock at the output of the MMCM. 
signal RESET: std_logic:='0'; -- Internal RESET after the clocks are stable  
signal USER_RESET: std_logic:='0'; -- User-controlled global reset
signal ALL_RESET: std_logic:='0'; -- Combined hard and soft global reset
signal SYSMON_CLK:   std_logic;
signal clk125_reset_reg: std_logic;

signal local_mac_addr: std_logic_vector(47 downto 0);
signal local_subarray: std_logic_vector(1 downto 0);
signal local_ip_addr: std_logic_vector(31 downto 0);
signal local_base_ip_port: std_logic_vector(15 downto 0);
signal remote_ip_port0: std_logic_vector(15 downto 0);
signal remote_ip_port1: std_logic_vector(15 downto 0);
-- Ethernet/UDP output / MASTER input  interface buses
signal axis_udp_tx_tdata:   std_logic_vector(7 downto 0);
signal axis_udp_tx_tlast:   std_logic;
signal axis_udp_tx_tvalid:   std_logic;
signal axis_udp_tx_tready:   std_logic;
signal udp0_tx_port:   std_logic_vector(1 downto 0) := (others=>'0');

signal axis_udp_rx_tdata: std_logic_vector(7 downto 0);
signal axis_udp_rx_tvalid: std_logic;
signal axis_udp_rx_tlast: std_logic;
signal axis_udp_rx_tready: std_logic;

signal sfp_tx_p: std_logic;
signal sfp_tx_n: std_logic;
signal sfp_rx_p: std_logic;
signal sfp_rx_n: std_logic;
signal sfp_refclk_nobuf: std_logic;
signal sfp_refclk_buf: std_logic;
signal sfp_status_vector_int: std_logic_vector(15 downto 0); -- Core status.
signal sfp_mmcm_locked: std_logic;
signal sfp_reset_done: std_logic;
signal udp_tx_overflow: std_logic;
signal udp_rx_overflow: std_logic;

signal lfsr_1 :std_logic_vector(7 downto 0);
signal lfsr_2 :std_logic_vector(7 downto 0);
----------------------------------------------------------------------------------
-- SYSTEM CLOCK
----------------------------------------------------------------------------------


component CLOCKS_V6 is
    PORT(
    -- Clock input
        SYSCLK_P : IN std_logic;
        SYSCLK_N : IN std_logic;

        
    -- General system clocks
        CLK25 : OUT std_logic;
        CLK200 : OUT std_logic;
        CLK200_MMCM_NOBUF : OUT std_logic; --! 200 MHz clock generated by a MMCM, *without* a BUFG. Is meant to be connected to the BUFGMUX that select the antenna processing clock. Cannot clock logic.
        CORR_CLK : OUT std_logic;
        PROC_CLK : OUT std_logic;
        CLK125 : OUT std_logic;
        SYSMON_CLK: OUT  STD_LOGIC; --! System monitor clock. Clocks the SYSMON hardware block. 

    -- Reset
        RST_IN : IN std_logic;          
        RST_OUT: OUT STD_LOGIC -- active high when everything is finished resseting
        );
end component;


component demo_funcgen is
    Port ( 
    --ce: in std_logic := '1'; 
    clk: in std_logic; -- clock period = 5.0 ns (200.0 Mhz)
    led: out std_logic_vector(7 downto 0)
    );
end component;


component hw7_3 is
  port (
    fir_in : in std_logic_vector( 8-1 downto 0 );
    clk : in std_logic;
    fir_out : out std_logic_vector( 8-1 downto 0 )
  );
end component;

component hw5_1_struct is
  port (
    gateway_in : in std_logic_vector( 16-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    gateway_out : out std_logic_vector( 8-1 downto 0 );
    gateway_out1 : out std_logic_vector( 8-1 downto 0 )
  );
end component;

  signal word_counter: unsigned(7 downto 0):=(others=>'0');
  signal ctr: unsigned(15 downto 0):=(others=>'0');-- X"00", to_unsigned(0,16)
  signal startup_ctr: unsigned(31 downto 0):=(others=>'0');
  signal wait_ctr: unsigned(15 downto 0):=(others=>'0');

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------


begin

--demo_funcgen0: demo_funcgen
--    port map(
     
--     clk => CLK125,
--     led => axis_udp_tx_tdata
     
--     );
     
     
hw5_uut: hw5_1_struct
  port map(
    gateway_in => "0000000000000000", --inital seed if you need to set it
    clk_1 => CLK125,
    ce_1 => '1',
    gateway_out => lfsr_1,
    gateway_out1 => lfsr_2
  );


hw7_uut: hw7_3 
  port map (
    fir_in => lfsr_1,
    clk => CLK125,
    fir_out => axis_udp_tx_tdata
  );


axis_udp_tx_tvalid<='1';
axis_udp_rx_tready<='1';
all_reset <= '0';
udp0_tx_port <= "00";
clk125_reset_reg <= '0';


  txproc: process(clk125)
  begin
    if rising_edge(clk125) then

      --if startup_ctr(31)='0' then
      --  startup_ctr<=startup_ctr+1;
      --  axis_udp_tx_tvalid<='0';
      --  axis_udp_rx_tready<='1';
      --else
        --if signed(wait_ctr(7 downto 0)) = 0 then -- 9 worked
            ctr<=ctr+1;

            --axis_udp_tx_tdata<=std_logic_vector(ctr(7 downto 0));
            if signed(ctr(10 downto 0))=-1 then
                axis_udp_tx_tlast<='1';
                --word_counter<=word_counter+1;
                --wait_ctr<=wait_ctr+1;
                GPIO_LED <= axis_udp_tx_tdata;
            else
                axis_udp_tx_tlast<='0';
            end if;                 
        --else
        --  wait_ctr<=wait_ctr+1;
        --  axis_udp_tx_tvalid<='0';
        --  axis_udp_rx_tready<='1';
        --end if;
      --end if;
     end if; --clk
  end process; 


--! Instantiate the system clock generator tht generates the local 200 MHz and 125 MHz from the external 200 MHz lines 
CLK0: CLOCKS_V6
    port map
        (
        -- System clock input
        SYSCLK_P=>SYSCLK_P,
        SYSCLK_N=>SYSCLK_N,
        -- Clocks using the internal clock manager
        CLK125 => CLK125,
        CLK200 => CLK200,
        CLK200_MMCM_NOBUF=>CLK200_MMCM_NOBUF,
        CLK25 => CLK25, -- generate 25 MHz clock for FMC board PLL reference
        CORR_CLK => CORR_CLK, -- Correlator clock
        SYSMON_CLK => SYSMON_CLK,
        
        -- Reset
        RST_IN=>ALL_RESET,
        RST_OUT=>RESET
        );





---------------------------------------------------------------------
-- UDP Interface on Marvell PHY
---------------------------------------------------------------------
--! Instantiate UDP / IP / Ethernet interface on PHY (Marvell Alaska) port
--! Keep to make sure the corresponding clocking ressources are used
local_mac_addr <= std_logic_vector'(X"12_34_56_78_9a_bc");


    udp_mac0: entity work.udp_mac
        GENERIC MAP(
            PHY_TYPE=> "GMII",  -- "GMII": Alaska 881111 PHY,  or "SGMII": SFP module
            SGMII_CLOCK_SOURCE => "0",  --SGMII_CLOCK_SOURCE,
            BROADCAST_IP_PORT => 41000, -- port on which broadcast requests and replies are made. This is fixed as it is used to discover the boards on the network and configure them.
            SIM => FALSE
            )
        PORT MAP(
            local_mac_addr =>local_mac_addr,
            local_ip_addr  =>X"0A0A0A0A",
            local_ip_port  =>X"A028",
            local_subarray => "00",
            -- User-side streaming interface
            remote_mac_addr =>X"0C4DE9A06A7A", -- Auto detect
            remote_ip_addr  =>X"0A0A0A0F", -- Auto detect
            remote_ip_port0  => X"A028", --remote_ip_port0, -- reply to port from the last incoming packet
            remote_ip_port1  => X"A029", --remote_ip_port1, -- reply to port from the last incoming packet

            -- GMII Phy interface (connects to Marvell chip pins)
            phy_rxclk        => phy_rxclk,
            phy_txer         => phy_txer,
            phy_reset_l      => phy_reset_l,
            phy_rxctrl_rxdv  => phy_rxctrl_rxdv,
            phy_rxd          => phy_rxd,
            phy_txc_gtxclk   => phy_txc_gtxclk, -- TX bus clock povided by the FPGA to the PHY
            phy_txctl_txen   => phy_txctl_txen,
            phy_txd          => phy_txd,
            phy_txclk        => phy_txclk, -- TX bus Clock provided *BY* the PHY for MII interfaces only. Not used.

            -- SGMII PHY interface (connects to SFP module pins and refernence clock source)
            -- sfp_clk_p => sfp_clk_p,
            -- sfp_clk_n => sfp_clk_n,
            sfp_tx_p => sfp_tx_p,
            sfp_tx_n => sfp_tx_n,
            sfp_rx_p => sfp_rx_p,
            sfp_rx_n => sfp_rx_n,

            -- SGMII buffered reference clock
            sfp_refclk_nobuf => sfp_refclk_nobuf, -- Unbuffered 125 MHz clock from the SFP reference clock.
            sfp_refclk_buf => sfp_refclk_buf, -- Buffered 125 MHz clock from the SFP reference clock.

            -- SGMII-specific status signals
            status_vector => sfp_status_vector_int,
            mmcm_locked => sfp_mmcm_locked,
            reset_done => sfp_reset_done,

            -- User TX interface
            s_axis_udp_tx_tvalid => axis_udp_tx_tvalid,
            s_axis_udp_tx_tdata  => axis_udp_tx_tdata,
            s_axis_udp_tx_tlast  => axis_udp_tx_tlast,
            s_axis_udp_tx_tready => axis_udp_tx_tready,
            tx_port              => udp0_tx_port,

            m_axis_udp_rx_tdata  => axis_udp_rx_tdata,
            m_axis_udp_rx_tvalid => axis_udp_rx_tvalid,
            m_axis_udp_rx_tlast  => axis_udp_rx_tlast,
            m_axis_udp_rx_tready => axis_udp_rx_tready,

            tx_overflow          => udp_tx_overflow,
            rx_overflow          => udp_rx_overflow,

            clk125 => clk125, -- User RX/TX interface clock AND GMII transmit clock (SGMII uses either this or th SFP reference clock). For SGMII, this must be a stable clock not related to any of the SGMII clocks.
            -- clk200 => clk200, -- used for the SGMII interface to initialize the cores even if the transceiver is not locked

            -- rst => ctrl_rst
            rst => clk125_reset_reg
        );


end Behavioral;

